library ieee;
  use ieee.std_logic_1164.all;




architecture scratch of led4_button4 is

  constant button_tab_c : natural := 1;



begin

  process(clk)
  begin
    if rising_edge(clk) then
      if reset = '1' then
        leds <= "0000";
      else
        leds() <= and(buttons);
        leds() <= or(buttons);
        leds() <= xor(buttons);
        leds() <= nor(buttons);
      end if;
    end if;
  end process;

end architecture;
