architecture scratch of led4_button4 is
begin
end architecture;
