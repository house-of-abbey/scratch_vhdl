-------------------------------------------------------------------------------------
--
-- Distributed under MIT Licence
--   See https://github.com/house-of-abbey/scratch_vhdl/blob/main/LICENCE.
--
-------------------------------------------------------------------------------------
--
-- This file is overwritten by Scratch VHDL code generation. We just need a stub in
-- order to add the file to a Vivado project.
--
-- J D Abbey & P A Abbey, 27 October 2022
--
-------------------------------------------------------------------------------------

architecture scratch of led4_button4 is
begin
end architecture;
