-------------------------------------------------------------------------------------
--
-- Distributed under MIT Licence
--   See https://github.com/house-of-abbey/scratch_vhdl/blob/main/LICENCE.
--
-------------------------------------------------------------------------------------
--
-- An empty scratch architecture solely for Vivado. This is deliberately excluded
-- from the ModelSim compilation.
--
-- J D Abbey & P A Abbey, 27 October 2022
--
-------------------------------------------------------------------------------------

architecture scratch of led4_button4 is
begin

  assert false
    report "Empty scratch architecture"
    severity failure;

end architecture;
